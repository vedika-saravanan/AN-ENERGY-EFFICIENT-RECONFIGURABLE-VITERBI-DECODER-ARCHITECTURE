library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all;
    
    
   entity sub is 
    
      port (
      
             in1 : in std_logic_vector ( 7 downto 0 ) ;
             in2 : in std_logic_vector ( 7 downto 0 ) ;               
             output : out std_logic_vector ( 8 downto 0 ) 
             
        ) ;
        
   end sub ;


architecture behav of sub is 

   begin       
       
        output <= ('0' & in1) - ('0' & in2) ;
        
end behav ;